module EnemyFleet
    (
    clk,
    reset,
    start,
    
    )